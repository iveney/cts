* spice from s1s
.include tuned_45nm_HP.pm
.subckt inv in out vdd
m1  out in  vdd vdd   pmos l=45n w=14.6u
m2  out in  0   0     nmos l=45n w=10.0u 
.ends inv
c0 n0 0 38.8889f
c1 n8 0 38.8888f
c2 n9 0 38.889f
c3 n10 0 38.8887f
c4 n11 0 38.8889f
c5 n12 0 38.8888f
c6 n13 0 42.5148f
c7 n1 0 105.8088f
c8 n14 0 31.6372f
c9 n15 0 37.7778f
c10 n16 0 31.6569f
c11 n17 0 34.4576f
c12 n2 0 44.4444f
c13 n22 0 3.3333f
c14 n23 0 38.8889f
c15 n24 0 3.3333f
c16 n25 0 38.8889f
c17 n5 0 61.0848f
c18 n18 0 13.3138f
c19 n19 0 38.8954f
c20 n20 0 13.3137f
c21 n21 0 38.8955f
c22 n3 0 73.8889f
c23 n4 0 73.8889f
c24 n6 0 73.8954f
c25 n7 0 73.8953f
c26 nSEG_NODE_26 0 77.7778f
c27 nSEG_NODE_27 0 77.7777f
c28 nSEG_NODE_28 0 77.778f
c29 nSEG_NODE_29 0 77.7777f
c30 nSEG_NODE_30 0 77.7778f
c31 nSEG_NODE_31 0 77.7777f
c32 nSEG_NODE_32 0 85.0295f
c33 nSEG_NODE_33 0 75.5556f
c34 nSEG_NODE_34 0 75.5556f
c35 nSEG_NODE_35 0 68.9152f
c36 nSEG_NODE_36 0 68.9149f
c37 nSEG_NODE_37 0 77.7778f
c38 nSEG_NODE_38 0 77.7778f
c39 nSEG_NODE_39 0 77.7778f
c40 nSEG_NODE_40 0 77.7778f
c41 nSEG_NODE_41 0 77.7908f
c42 nSEG_NODE_42 0 77.7908f
c43 nSEG_NODE_43 0 77.791f
c44 nSEG_NODE_44 0 77.7908f
r0 n0 n8 116.6666
r1 n9 n10 116.6667
r2 n11 n12 116.6666
r3 n13 n1 85.0295
r4 n1 n14 31.6372
r5 n15 n2 113.3334
r6 n1 n16 31.6569
r7 n17 n5 103.3725
r8 n2 n22 3.3333
r9 n23 n3 116.6667
r10 n2 n24 3.3333
r11 n25 n4 116.6667
r12 n5 n18 13.3138
r13 n19 n6 116.6862
r14 n5 n20 13.3137
r15 n21 n7 116.6863
r16 n0 nSEG_NODE_26 38.8889
r17 nSEG_NODE_26 nSEG_NODE_27 38.8889
r18 nSEG_NODE_27 n8 38.8888
r19 n9 nSEG_NODE_28 38.889
r20 nSEG_NODE_28 nSEG_NODE_29 38.889
r21 nSEG_NODE_29 n10 38.8887
r22 n11 nSEG_NODE_30 38.8889
r23 nSEG_NODE_30 nSEG_NODE_31 38.8889
r24 nSEG_NODE_31 n12 38.8888
r25 n13 nSEG_NODE_32 42.5148
r26 nSEG_NODE_32 n1 42.5147
r27 n15 nSEG_NODE_33 37.7778
r28 nSEG_NODE_33 nSEG_NODE_34 37.7778
r29 nSEG_NODE_34 n2 37.7778
r30 n17 nSEG_NODE_35 34.4576
r31 nSEG_NODE_35 nSEG_NODE_36 34.4576
r32 nSEG_NODE_36 n5 34.4573
r33 n23 nSEG_NODE_37 38.8889
r34 nSEG_NODE_37 nSEG_NODE_38 38.8889
r35 nSEG_NODE_38 n3 38.8889
r36 n25 nSEG_NODE_39 38.8889
r37 nSEG_NODE_39 nSEG_NODE_40 38.8889
r38 nSEG_NODE_40 n4 38.8889
r39 n19 nSEG_NODE_41 38.8954
r40 nSEG_NODE_41 nSEG_NODE_42 38.8954
r41 nSEG_NODE_42 n6 38.8954
r42 n21 nSEG_NODE_43 38.8955
r43 nSEG_NODE_43 nSEG_NODE_44 38.8955
r44 nSEG_NODE_44 n7 38.8953
x0 gin n0 vdd inv
x1 n8 n9 vdd inv
x2 n10 n11 vdd inv
x3 n12 n13 vdd inv
x4 n14 n15 vdd inv
x5 n22 n23 vdd inv
x6 n24 n25 vdd inv
x7 n16 n17 vdd inv
x8 n18 n19 vdd inv
x9 n20 n21 vdd inv
*
vdd vdd 0 1
vdt gin 0 1 pwl(0n 1, 0.2n 1, 0.325n 0, 2n 0)
*
.ic v(gin)=1
.ic v(n0)=0
.ic v(n8)=0
.ic v(n9)=1
.ic v(n10)=1
.ic v(n11)=0
.ic v(n12)=0
.ic v(n13)=1
.ic v(n1)=1
.ic v(n14)=1
.ic v(n15)=0
.ic v(n16)=1
.ic v(n17)=0
.ic v(n2)=0
.ic v(n22)=0
.ic v(n23)=1
.ic v(n24)=0
.ic v(n25)=1
.ic v(n5)=0
.ic v(n18)=0
.ic v(n19)=1
.ic v(n20)=0
.ic v(n21)=1
.ic v(n3)=1
.ic v(n4)=1
.ic v(n6)=1
.ic v(n7)=1
.ic v(nSEG_NODE_26)=0
.ic v(nSEG_NODE_27)=0
.ic v(nSEG_NODE_28)=0
.ic v(nSEG_NODE_29)=0
.ic v(nSEG_NODE_30)=0
.ic v(nSEG_NODE_31)=0
.ic v(nSEG_NODE_32)=0
.ic v(nSEG_NODE_33)=0
.ic v(nSEG_NODE_34)=0
.ic v(nSEG_NODE_35)=0
.ic v(nSEG_NODE_36)=0
.ic v(nSEG_NODE_37)=0
.ic v(nSEG_NODE_38)=0
.ic v(nSEG_NODE_39)=0
.ic v(nSEG_NODE_40)=0
.ic v(nSEG_NODE_41)=0
.ic v(nSEG_NODE_42)=0
.ic v(nSEG_NODE_43)=0
.ic v(nSEG_NODE_44)=0
*
.opti nopage temp=75
.width out=240
*
.tran 0.01n 2n 0.0n 0.01n
.print tran v(gin) v(n8) v(n10) v(n12) v(n14) v(n22) v(n24) v(n16) v(n18) v(n20) v(n3) v(n4) v(n6) v(n7)
* plot v(gin) v(n8) v(n10) v(n12) v(n14) v(n22) v(n24) v(n16) v(n18) v(n20) v(n3) v(n4) v(n6) v(n7)
.end
