* spice from s2s
.include tuned_45nm_HP.pm
.subckt inv in out vdd
m1  out in  vdd vdd   pmos l=45n w=14.6u
m2  out in  0   0     nmos l=45n w=10.0u 
.ends inv
c0 n0 0 36.6313f
c1 n16 0 36.6313f
c2 n17 0 36.6314f
c3 n18 0 36.6313f
c4 n19 0 36.6314f
c5 n20 0 36.6313f
c6 n21 0 36.6313f
c7 n22 0 36.6313f
c8 n23 0 36.6314f
c9 n24 0 36.6313f
c10 n25 0 36.6314f
c11 n26 0 36.6313f
c12 n27 0 36.6314f
c13 n28 0 36.6313f
c14 n29 0 28.6459f
c15 n1 0 64.9649f
c16 n34 0 26.6378f
c17 n35 0 36.8559f
c18 n36 0 36.8556f
c19 n37 0 36.8558f
c20 n50 0 36.8558f
c21 n51 0 36.8558f
c22 n52 0 36.8558f
c23 n53 0 36.8558f
c24 n3 0 46.4301f
c25 n32 0 30.4592f
c26 n33 0 48.7162f
c27 n38 0 48.7161f
c28 n39 0 48.7162f
c29 n48 0 48.7161f
c30 n49 0 48.7161f
c31 n54 0 48.7161f
c32 n55 0 28.7162f
c33 n30 0 6.2896f
c34 n31 0 28.0015f
c35 n4 0 108.7161f
c36 n7 0 70.1387f
c37 n40 0 17.2597f
c38 n41 0 36.6314f
c39 n46 0 36.6313f
c40 n47 0 39.242f
c41 n42 0 24.8775f
c42 n43 0 40.4403f
c43 n44 0 40.4403f
c44 n45 0 31.761f
c45 n8 0 120.0001f
c46 n58 0 46.7373f
c47 n59 0 42.9896f
c48 n56 0 34.0208f
c49 n57 0 48.2627f
c50 n10 0 98.2627f
c51 n13 0 129.9999f
c52 n60 0 49.1195f
c53 n61 0 40.4403f
c54 n62 0 49.1194f
c55 n63 0 40.4403f
c56 n2 0 71.8558f
c57 n5 0 75f
c58 n6 0 75f
c59 n9 0 77.9896f
c60 n11 0 60f
c61 n12 0 60f
c62 n14 0 75.4402f
c63 n15 0 75.4403f
c64 nSEG_NODE_64 0 73.2626f
c65 nSEG_NODE_65 0 73.2627f
c66 nSEG_NODE_66 0 73.2627f
c67 nSEG_NODE_67 0 73.2626f
c68 nSEG_NODE_68 0 73.2627f
c69 nSEG_NODE_69 0 73.2627f
c70 nSEG_NODE_70 0 73.2627f
c71 nSEG_NODE_71 0 57.2917f
c72 nSEG_NODE_72 0 53.2756f
c73 nSEG_NODE_73 0 73.7118f
c74 nSEG_NODE_74 0 73.7115f
c75 nSEG_NODE_75 0 73.7116f
c76 nSEG_NODE_76 0 73.7116f
c77 nSEG_NODE_77 0 73.7116f
c78 nSEG_NODE_78 0 73.7116f
c79 nSEG_NODE_79 0 73.7116f
c80 nSEG_NODE_80 0 73.7116f
c81 nSEG_NODE_81 0 97.4323f
c82 nSEG_NODE_82 0 97.4323f
c83 nSEG_NODE_83 0 97.4322f
c84 nSEG_NODE_84 0 57.4323f
c85 nSEG_NODE_85 0 56.003f
c86 nSEG_NODE_86 0 73.2627f
c87 nSEG_NODE_87 0 80.8806f
c88 nSEG_NODE_88 0 85.9792f
c89 nSEG_NODE_89 0 80.8805f
c90 nSEG_NODE_90 0 80.8806f
r0 n0 n16 73.2626
r1 n17 n18 73.2627
r2 n19 n20 73.2627
r3 n21 n22 73.2626
r4 n23 n24 73.2627
r5 n25 n26 73.2627
r6 n27 n28 73.2627
r7 n29 n1 57.2917
r8 n1 n34 53.2756
r9 n35 n36 110.5674
r10 n37 n50 110.5674
r11 n51 n52 110.5674
r12 n53 n2 110.5674
r13 n1 n3 9.6813
r14 n3 n32 30.4592
r15 n33 n38 97.4323
r16 n39 n48 97.4323
r17 n49 n54 97.4322
r18 n55 n4 57.4323
r19 n3 n30 6.2896
r20 n31 n7 56.003
r21 n4 n5 40
r22 n4 n6 40
r23 n7 n40 17.2597
r24 n41 n46 73.2627
r25 n47 n8 39.242
r26 n7 n42 24.8775
r27 n43 n44 80.8806
r28 n45 n13 31.761
r29 n8 n58 46.7373
r30 n59 n9 85.9792
r31 n8 n56 34.0208
r32 n57 n10 48.2627
r33 n10 n11 25
r34 n10 n12 25
r35 n13 n60 49.1195
r36 n61 n14 80.8805
r37 n13 n62 49.1194
r38 n63 n15 80.8806
r39 n0 nSEG_NODE_64 36.6313
r40 nSEG_NODE_64 n16 36.6313
r41 n17 nSEG_NODE_65 36.6314
r42 nSEG_NODE_65 n18 36.6313
r43 n19 nSEG_NODE_66 36.6314
r44 nSEG_NODE_66 n20 36.6313
r45 n21 nSEG_NODE_67 36.6313
r46 nSEG_NODE_67 n22 36.6313
r47 n23 nSEG_NODE_68 36.6314
r48 nSEG_NODE_68 n24 36.6313
r49 n25 nSEG_NODE_69 36.6314
r50 nSEG_NODE_69 n26 36.6313
r51 n27 nSEG_NODE_70 36.6314
r52 nSEG_NODE_70 n28 36.6313
r53 n29 nSEG_NODE_71 28.6459
r54 nSEG_NODE_71 n1 28.6458
r55 n1 nSEG_NODE_72 26.6378
r56 nSEG_NODE_72 n34 26.6378
r57 n35 nSEG_NODE_73 36.8559
r58 nSEG_NODE_73 nSEG_NODE_74 36.8559
r59 nSEG_NODE_74 n36 36.8556
r60 n37 nSEG_NODE_75 36.8558
r61 nSEG_NODE_75 nSEG_NODE_76 36.8558
r62 nSEG_NODE_76 n50 36.8558
r63 n51 nSEG_NODE_77 36.8558
r64 nSEG_NODE_77 nSEG_NODE_78 36.8558
r65 nSEG_NODE_78 n52 36.8558
r66 n53 nSEG_NODE_79 36.8558
r67 nSEG_NODE_79 nSEG_NODE_80 36.8558
r68 nSEG_NODE_80 n2 36.8558
r69 n33 nSEG_NODE_81 48.7162
r70 nSEG_NODE_81 n38 48.7161
r71 n39 nSEG_NODE_82 48.7162
r72 nSEG_NODE_82 n48 48.7161
r73 n49 nSEG_NODE_83 48.7161
r74 nSEG_NODE_83 n54 48.7161
r75 n55 nSEG_NODE_84 28.7162
r76 nSEG_NODE_84 n4 28.7161
r77 n31 nSEG_NODE_85 28.0015
r78 nSEG_NODE_85 n7 28.0015
r79 n41 nSEG_NODE_86 36.6314
r80 nSEG_NODE_86 n46 36.6313
r81 n43 nSEG_NODE_87 40.4403
r82 nSEG_NODE_87 n44 40.4403
r83 n59 nSEG_NODE_88 42.9896
r84 nSEG_NODE_88 n9 42.9896
r85 n61 nSEG_NODE_89 40.4403
r86 nSEG_NODE_89 n14 40.4402
r87 n63 nSEG_NODE_90 40.4403
r88 nSEG_NODE_90 n15 40.4403
x0 gin n0 vdd inv
x1 n16 n17 vdd inv
x2 n18 n19 vdd inv
x3 n20 n21 vdd inv
x4 n22 n23 vdd inv
x5 n24 n25 vdd inv
x6 n26 n27 vdd inv
x7 n28 n29 vdd inv
x8 n28 n29 vdd inv
x9 n34 n35 vdd inv
x10 n36 n37 vdd inv
x11 n50 n51 vdd inv
x12 n52 n53 vdd inv
x13 n52 n53 vdd inv
x14 n32 n33 vdd inv
x15 n38 n39 vdd inv
x16 n48 n49 vdd inv
x17 n54 n55 vdd inv
x18 n54 n55 vdd inv
x19 n30 n31 vdd inv
x20 n30 n31 vdd inv
x21 n40 n41 vdd inv
x22 n46 n47 vdd inv
x23 n46 n47 vdd inv
x24 n58 n59 vdd inv
x25 n58 n59 vdd inv
x26 n56 n57 vdd inv
x27 n56 n57 vdd inv
x28 n42 n43 vdd inv
x29 n44 n45 vdd inv
x30 n44 n45 vdd inv
x31 n60 n61 vdd inv
x32 n60 n61 vdd inv
x33 n62 n63 vdd inv
x34 n62 n63 vdd inv
*
vdd vdd 0 1.2
vdt gin 0 1.2 pwl(0n 1.2, 0.2n 1.2, 0.325n 0, 2n 0)
*
.ic v(gin)=1.2
.ic v(n0)=0
.ic v(n16)=0
.ic v(n17)=1.2
.ic v(n18)=1.2
.ic v(n19)=0
.ic v(n20)=0
.ic v(n21)=1.2
.ic v(n22)=1.2
.ic v(n23)=0
.ic v(n24)=0
.ic v(n25)=1.2
.ic v(n26)=1.2
.ic v(n27)=0
.ic v(n28)=0
.ic v(n29)=1.2
.ic v(n1)=1.2
.ic v(n34)=1.2
.ic v(n35)=0
.ic v(n36)=0
.ic v(n37)=1.2
.ic v(n50)=1.2
.ic v(n51)=0
.ic v(n52)=0
.ic v(n53)=1.2
.ic v(n3)=1.2
.ic v(n32)=1.2
.ic v(n33)=0
.ic v(n38)=0
.ic v(n39)=1.2
.ic v(n48)=1.2
.ic v(n49)=0
.ic v(n54)=0
.ic v(n55)=1.2
.ic v(n30)=1.2
.ic v(n31)=0
.ic v(n4)=1.2
.ic v(n7)=0
.ic v(n40)=0
.ic v(n41)=1.2
.ic v(n46)=1.2
.ic v(n47)=0
.ic v(n42)=0
.ic v(n43)=1.2
.ic v(n44)=1.2
.ic v(n45)=0
.ic v(n8)=0
.ic v(n58)=0
.ic v(n59)=1.2
.ic v(n56)=0
.ic v(n57)=1.2
.ic v(n10)=1.2
.ic v(n13)=0
.ic v(n60)=0
.ic v(n61)=1.2
.ic v(n62)=0
.ic v(n63)=1.2
.ic v(n2)=1.2
.ic v(n5)=1.2
.ic v(n6)=1.2
.ic v(n9)=1.2
.ic v(n11)=1.2
.ic v(n12)=1.2
.ic v(n14)=1.2
.ic v(n15)=1.2
.ic v(nSEG_NODE_64)=0
.ic v(nSEG_NODE_65)=0
.ic v(nSEG_NODE_66)=0
.ic v(nSEG_NODE_67)=0
.ic v(nSEG_NODE_68)=0
.ic v(nSEG_NODE_69)=0
.ic v(nSEG_NODE_70)=0
.ic v(nSEG_NODE_71)=0
.ic v(nSEG_NODE_72)=0
.ic v(nSEG_NODE_73)=0
.ic v(nSEG_NODE_74)=0
.ic v(nSEG_NODE_75)=0
.ic v(nSEG_NODE_76)=0
.ic v(nSEG_NODE_77)=0
.ic v(nSEG_NODE_78)=0
.ic v(nSEG_NODE_79)=0
.ic v(nSEG_NODE_80)=0
.ic v(nSEG_NODE_81)=0
.ic v(nSEG_NODE_82)=0
.ic v(nSEG_NODE_83)=0
.ic v(nSEG_NODE_84)=0
.ic v(nSEG_NODE_85)=0
.ic v(nSEG_NODE_86)=0
.ic v(nSEG_NODE_87)=0
.ic v(nSEG_NODE_88)=0
.ic v(nSEG_NODE_89)=0
.ic v(nSEG_NODE_90)=0
*
.opti nopage temp=75
.width out=240
*
.tran 0.01n 2n 0.0n 0.01n
.print tran v(gin) v(n16) v(n18) v(n20) v(n22) v(n24) v(n26) v(n28) v(n34) v(n36) v(n50) v(n52) v(n32) v(n38) v(n48) v(n54) v(n30) v(n40) v(n46) v(n58) v(n56) v(n42) v(n44) v(n60) v(n62) v(n2) v(n5) v(n6) v(n9) v(n11) v(n12) v(n14) v(n15)
* plot v(gin) v(n16) v(n18) v(n20) v(n22) v(n24) v(n26) v(n28) v(n34) v(n36) v(n50) v(n52) v(n32) v(n38) v(n48) v(n54) v(n30) v(n40) v(n46) v(n58) v(n56) v(n42) v(n44) v(n60) v(n62) v(n2) v(n5) v(n6) v(n9) v(n11) v(n12) v(n14) v(n15)
.end
